//XOR Gate
//Structural modelling

module XOR_Structural(a,b,y);
input a,b;
output y;

xor xor1(y,a,b);
endmodule
