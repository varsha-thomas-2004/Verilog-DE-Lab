//OR Gate
//Structural modelling

module OR_Structural(a,b,y);
input a,b;
output y;

or or1(y,a,b);

endmodule
