//NOT Gate
//Structural modelling

module NOT_Structural(a,y);
input a;
output y;

not not1(y,a);

endmodule
