//NOT Gate
//Dataflow modelling

module NOT_Dataflow(a,y);
input a;
output y;

assign y = ~a;
endmodule
