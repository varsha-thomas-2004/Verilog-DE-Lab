//AND Gate
//Dataflow modelling

module AND_Dataflow(a,b,y);
input a,b;
output y;

assign y = a & b;

endmodule
