//AND Gate
//Structural modelling

module AND(a,b,y);
input a,b;
output y;

and and1(y,a,b);

endmodule 